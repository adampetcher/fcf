(* Copyright 2012-2015 by Adam Petcher.				*
 * Use of this source code is governed by the license described	*
 * in the LICENSE file at the root of the source tree.		*)
(* A top-level module that exports all of the common components of the framework. *)

Require Export FCF.DistRules.
Require Export FCF.Comp.
Require Export Arith.
Require Export FCF.Fold.
Require Export FCF.Rat.
Require Export FCF.DistSem.
Require Export FCF.StdNat.
Require Export FCF.DistTacs.


Open Scope comp_scope.
Open Scope rat_scope.
