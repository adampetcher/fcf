(* Copyright 2012-2015 by Adam Petcher.				*
 * Use of this source code is governed by the license described	*
 * in the LICENSE file at the root of the source tree.		*)
(* A top-level module that exports all of the common components of the framework. *)

Require Export DistRules.
Require Export Comp.
Require Export Arith.
Require Export Fold.
Require Export Rat.
Require Export DistSem.
Require Export StdNat.
Require Export DistTacs.


Open Scope comp_scope.
Open Scope rat_scope.